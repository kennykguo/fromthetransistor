module hello; initial $display ("Hello World!"); endmodule
./obj_dir/Vhello